//-----------------------------------------------------
// File Name   : alucodes.sv
// Function    : pMIPS ALU function code definitions 
// Author:   tjk
// Last rev. 23 Oct 12 
//-----------------------------------------------------
// 
`define RADD  3'b010
`define RSUB  3'b011  
`define RMUL 3'b100